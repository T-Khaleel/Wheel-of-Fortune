library verilog;
use verilog.vl_types.all;
entity wof_vlg_vec_tst is
end wof_vlg_vec_tst;
